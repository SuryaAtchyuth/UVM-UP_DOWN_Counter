
interface count_interface(input clk);

  logic      rst;
  logic[3:0] out;
  
endinterface: count_interface  
  
